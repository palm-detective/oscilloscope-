* model for lmh6643max
* see orginal LMH6643 model from National Semi
* PAA 08/2021
**********************************************************
.OPTIONS  ACCT   LIST

.inc LMH6643.MOD
.subcircuit lmh6643max 1 2 3 4 5 6 7 8
LMH6643 2 3 8 4 1
LMH6643 6 5 8 4 7
.end

.ENDS
