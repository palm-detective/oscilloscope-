* model for HC4053
* Based on NXP models
* see notes for orginal NXP models
* PAA 05/2021
**********************************************************
.OPTIONS  ACCT   LIST

* Nominal parameters
.INC hc_tnomi.cir

* Fast parameters
*.INC hc_tfast.cir

* Slow parameters
*.INC hc_tslow.cir

**********************************************************
* Package Options
**********************************************************
*.INC ssop.s
*.INC so.s
*.INC dip.s
.INC tssop.s
*.INC dhvqfn.s

.SUBCKT HC4053 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
XHC4053A   40  50  60  70  80  90  SWI1
XHC4053B   41  51  61  70  80  90  SWI1
XHC4053C   42  52  62  70  80  90  SWI1
XPK16  1  2  3  4  5  6  7  0  9 10 11 12 13 14 15 16
+     51 61 62 42 52 20 70 90 90 90 90 50 60 40 41 80 pk16
* PIN  1  2  3  4  5  6  7  8  9 10 11 12 13 14 15 16
*     B1 B0 C1 CC C0  E V- GD SC SB SA A0 A1 AC BC V+
.ENDS

.end